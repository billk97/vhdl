library verilog;
use verilog.vl_types.all;
entity erg1_vlg_vec_tst is
end erg1_vlg_vec_tst;
