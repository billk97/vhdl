LIBRARY ieee;
USE ieee.std_logic_1164.all;
	ENTITY AXORB IS 
		PORT (MuxA,MuxB : IN STD_LOGIC;
				A_XOR_B : OUT STD_LOGIC );
		END AXORB;
	ARCHITECTURE ArchAXORB OF AXORB IS
		BEGIN 
			A_XOR_B  <=(MuxA AND (NOT MUXB))OR((NOT MUXA) AND MUXB);
		END ArchAXORB;