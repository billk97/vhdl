library verilog;
use verilog.vl_types.all;
entity erg3_vlg_vec_tst is
end erg3_vlg_vec_tst;
