library verilog;
use verilog.vl_types.all;
entity erg2_vlg_vec_tst is
end erg2_vlg_vec_tst;
